`define SIMMEM_DATA_WIDTH 64
`define MAX_NUM_LANES 32
`define SIMMEM_SOURCE_WIDTH 32
`define SIMMEM_LOGSIZE_WIDTH 8
